////////////////////////////////////////////////////////////////////////////////
// Module:  forward_unit.v
// Project: SJSU EE275 Mini Project 2
// Description: Forwarding control unit
//
// Name: Zach Smith 
// Student ID: 007159087
//
////////////////////////////////////////////////////////////////////////////////
`include "mips_defs.vh"

module forward_unit(
   
);

endmodule // forward_unit