////////////////////////////////////////////////////////////////////////////////
// File:  alu.vh
// Project: SJSU EE275 Mini Project 2
// Description:
//
// Name: Zach Smith 
// Student ID: 007159087
//
// Notes:
//
////////////////////////////////////////////////////////////////////////////////
`ifndef _ALU_VH
`define _ALU_VH

`define ALU_ADD   4'b0000
`define ALU_ADDU  4'b0001
`define ALU_SUB   4'b0010
`define ALU_SUBU  4'b0011
`define ALU_AND   4'b0100
`define ALU_OR    4'b0101
`define ALU_SLT   4'b0110
`define ALU_SLTU  4'b0111
`define ALU_FCN   4'b1000

`endif // _ALU_VH