////////////////////////////////////////////////////////////////////////////////
// Module:  mips_datapath.v
// Project: SJSU EE275 Mini Project 2
// Description: Portion of a 5-stage pipeline MIPS datapath with forwarding
//
// Name: Zach Smith 
// Student ID: 007159087
//
// Note:
//
////////////////////////////////////////////////////////////////////////////////

module mips_datapath(

);
parameter instruction_mem = "";
parameter data_mem = "";

endmodule // mips_datapath